:Address:City:Country:Employees:ID:Name:State:Latitude:Longitude:ZIP
0:3666 21st St:San Francisco:USA:8:1:Madeira:CA:37.756488877551:-122.429343346939:94114
1:735 Dolores St:San Francisco:USA:15:2:Bready Shop:CA:Unknown:Unknown:94119
2:332 Hill St:San Francisco:USA:25:3:Super River:California:37.755725122449:-122.428601306122:94114
3:3995 23rd St:San Francisco:USA:10:4:Ben's Shop:CA:37.7529648:-122.431714:94114
4:1056 Sanchez St:San Francisco:USA:12:5:Sanchez:California:37.7521458:-122.42981516:N/A
5:551 Alvarado St:San Francisco:USA:20:6:Richvalley:CA:37.7536733265306:-122.433219959184:94114
